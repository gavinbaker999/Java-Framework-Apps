entity test is
end test;
architecture testhdl of test is
end testhdl;
