entity ptest is
one: process(in1,in2)
end ptest;
