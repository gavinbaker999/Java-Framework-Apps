pOrt MAp if i++ (12.47) "this is a string" THen Q<='0';